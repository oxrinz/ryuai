module UART_TX (
    input            i_Rst_L,
    input            i_Clock,
    input            i_TX_DV,
    input      [7:0] i_TX_Byte,
    output reg       o_TX_Active,
    output reg       o_TX_Serial,
    output reg       o_TX_Done
);

  localparam IDLE = 2'b00;
  localparam TX_START_BIT = 2'b01;
  localparam TX_DATA_BITS = 2'b10;
  localparam TX_STOP_BIT = 2'b11;
  localparam CLKS_PER_BIT = 217;

  reg [2:0] r_SM_Main;
  reg [$clog2(CLKS_PER_BIT):0] r_Clock_Count;
  reg [2:0] r_Bit_Index;
  reg [7:0] r_TX_Data;

  always @(posedge i_Clock or negedge i_Rst_L) begin
    if (~i_Rst_L) begin
      r_SM_Main <= 3'b000;
    end else begin

      o_TX_Done <= 1'b0;

      case (r_SM_Main)
        IDLE: begin
          o_TX_Serial   <= 1'b1;
          r_Clock_Count <= 0;
          r_Bit_Index   <= 0;

          if (i_TX_DV == 1'b1) begin
            o_TX_Active <= 1'b1;
            r_TX_Data   <= i_TX_Byte;
            r_SM_Main   <= TX_START_BIT;
          end else r_SM_Main <= IDLE;
        end

        TX_START_BIT: begin
          o_TX_Serial <= 1'b0;

          if (r_Clock_Count < CLKS_PER_BIT - 1) begin
            r_Clock_Count <= r_Clock_Count + 1;
            r_SM_Main     <= TX_START_BIT;
          end else begin
            r_Clock_Count <= 0;
            r_SM_Main     <= TX_DATA_BITS;
          end
        end

        TX_DATA_BITS: begin
          o_TX_Serial <= r_TX_Data[r_Bit_Index];

          if (r_Clock_Count < CLKS_PER_BIT - 1) begin
            r_Clock_Count <= r_Clock_Count + 1;
            r_SM_Main     <= TX_DATA_BITS;
          end else begin
            r_Clock_Count <= 0;

            if (r_Bit_Index < 7) begin
              r_Bit_Index <= r_Bit_Index + 1;
              r_SM_Main   <= TX_DATA_BITS;
            end else begin
              r_Bit_Index <= 0;
              r_SM_Main   <= TX_STOP_BIT;
            end
          end
        end

        TX_STOP_BIT: begin
          o_TX_Serial <= 1'b1;

          if (r_Clock_Count < CLKS_PER_BIT - 1) begin
            r_Clock_Count <= r_Clock_Count + 1;
            r_SM_Main     <= TX_STOP_BIT;
          end else begin
            o_TX_Done     <= 1'b1;
            r_Clock_Count <= 0;
            r_SM_Main     <= IDLE;
            o_TX_Active   <= 1'b0;
          end
        end

        default: r_SM_Main <= IDLE;

      endcase
    end
  end

endmodule
