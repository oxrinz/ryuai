module PC ();



endmodule
